package yapp_pkg;
	import uvm_pkg::*;        //import UVM package
	`include "uvm_macros.svh" //include UVM macro file
	`include "yapp_packet.sv" //include design file
endpackage
